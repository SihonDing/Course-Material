library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Counter8 is
	port (clk: in std_logic;
	q: out std_logic_vector (2 downto 0)
	);
end Counter8;

architecture arch_Counter8 of Counter8 is
	signal tmp_q: std_logic_vector(2 downto 0) := "000";
begin
	q <= tmp_q;
	process(clk)
	begin
		if (clk'event and clk='1') then
			if (tmp_q="111") then
				tmp_q <= "000";
			else 
				tmp_q <= tmp_q + 1;
			end if;
		end if;
	end process;
end arch_Counter8;